`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 10/22/2023 02:05:28 PM
// Design Name: 
// Module Name: puf_challenge_response
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////

// -----------------------------------------------------------------------------
// Module: puf_challenge_response
//
// Description:
// This module implements a Finite State Machine (FSM) to interact with a 
// Physically Unclonable Function (PUF). The FSM takes a 6-bit challenge as 
// input and produces an 8-bit response based on the PUF's behavior. The FSM 
// transitions through several states including IDLE, START, WAIT, STORE, 
// INCREMENT, and COMPARE to manage the PUF operation and generate the response.
//
// Ports:
// - CLK: Clock input
// - recalculate: Signal to recalculate the response
// - challenge_lower_bits: Lower 6 bits of the challenge
// - response: 8-bit response generated by the FSM
// - completed: Signal to indicate completion of challenge-response
// -----------------------------------------------------------------------------

`define TRUE    1'b1
`define FALSE   1'b0
`define num_RO  8
// This is working. But does not help the PUF drifting problem.
// Modify the MAX_STD_COUNT in configurable_RO_PUF instead.
`define NUM_REPEAT 1   

module puf_challenge_response(
    input logic CLK,                    // Clock input
    input logic recalculate,            // Signal to recalculate the response
    input [5:0] challenge_lower_bits,   // Lower 6 bits of the challenge
    output logic [7:0] response,        // 8-bit response
    output logic completed              // Signal to indicate completion
);

    // Define FSM states
    typedef enum logic [3:0] {
        IDLE = 4'b0000,
        START,
        WAIT,
        STORE,
        INCREMENT,
        COMPARE
    } fsm_state_t;

    // Initialize current and next FSM states
    fsm_state_t state = IDLE, next_state;  
    
    // Declare and initialize internal signals and variables
    logic [31:0] ro_count_out;           // 32-bit counter output from PUF
    logic [9:0] challenge;               // 10-bit challenge input to PUF
    logic count_complete;                // Signal indicating PUF operation complete
    logic comparison_done;               // Flag for comparison completion
    logic [31:0] ro_count_array [8:0];   // Array to store ro_count_out values
    logic [3:0] index = 4'b0000;         // Index for array and upper 4 bits of challenge
    logic [5:0] prev_challenge_lower_bits; // Previous switch configuration
    logic [3:0] repeat_counter = 4'b0000;  // Counter for repetitions


    // FSM state transition logic
    always_ff @(posedge CLK) begin
        state <= next_state;
        prev_challenge_lower_bits <= challenge_lower_bits;  // Store current switch config for next cycle
    end

    // Next state logic based on current state and conditions
    always_comb begin
        next_state = state;
        case(state)
            IDLE:                           next_state = START;
            START:                          next_state = WAIT;
            WAIT:       if (count_complete) next_state = STORE;
            STORE:                          next_state = INCREMENT;
            INCREMENT:  if (index < `num_RO) next_state = START;
                        else                next_state = COMPARE;
            COMPARE:    if (comparison_done) begin
                            if ((prev_challenge_lower_bits != challenge_lower_bits) || recalculate) 
                                            next_state = IDLE;  // Transition to IDLE if switch config changed or recalculate is true
                            else
                                            next_state = COMPARE;  // Loop in COMPARE if switch config is the same
                        end
            default:    next_state = IDLE;
        endcase        
    end

    // Sequential Logic for FSM states
    always_ff @(posedge CLK) begin
        if (state == IDLE) begin
            index <= 4'b0000; // Reset upper challenges
            comparison_done <= `FALSE; // Reset flag at the beginning of each cycle
            
            
        end else if (state == START) begin
            challenge = {index, challenge_lower_bits}; // Update challenge bits
               
        end else if (state == STORE) begin            
            // Only average if the index will not increment
            if (repeat_counter < `NUM_REPEAT - 1) begin
                ro_count_array[index] <= (ro_count_out + ro_count_array[index]) >> 1;  
            end else begin
                ro_count_array[index] <= ro_count_out;
            end
            
            
        end else if (state == INCREMENT) begin
            if (repeat_counter >= `NUM_REPEAT - 1) begin
                index <= index + 1;  // Increment index for challenge bit
                repeat_counter <= 0;  // Reset the repeat counter
            end else begin
                repeat_counter <= repeat_counter + 1;  // Increment the repeat counter
            end
            
        end else if (state == COMPARE) begin // Compare counters and generate response
            for (int i = 0; i < `num_RO ; i = i + 1) begin
                response[i] <= (ro_count_array[i] < ro_count_array[i+1]) ? `TRUE : `FALSE;
            end            
            comparison_done <= `TRUE; // Set flag
        end
    end

    // Instantiate configurable_RO_PUF
    logic enable_ro_puf;  // Declare a new logic variable for the enable signal
    assign enable_ro_puf = (state != START) && (state != IDLE) && (state != COMPARE);
    configurable_RO_PUF puf_inst (
        .challenge(challenge),
        .clk(CLK),
        .en(enable_ro_puf),
        .ro_count_out(ro_count_out),
        .completed(count_complete)
    );
    
    // Assign the completed signal to indicate when challenge-response is done
    assign completed = comparison_done;
 
endmodule

